module hello();

	$display("hello world")

endmodule
